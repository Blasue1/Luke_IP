package simple_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "simple_trans.sv"
  `include "simple_sequence.sv"
  `include "simple_driver.sv"
  `include "simple_monitor.sv"
  `include "simple_scoreboard.sv"
  `include "simple_sequencer.sv"
  `include "simple_agent.sv"
  `include "simple_env.sv"
  `include "simple_test.sv"

endpackage
